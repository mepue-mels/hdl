module Testbench;
	initial begin 
		$display("Hi world");
	end
endmodule
